`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/04/2017 10:08:42 PM
// Design Name: 
// Module Name: RISC_V_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_RISC_V ;
// clock and reset signal declaration
    logic clk , reset ;
    logic [63:0] tb_ALU_Result ;
    logic  [31:0] INS_out;
    logic [63:0] mux_out;
    logic [63:0] rd1_out;
    logic [63:0] rd2_out;
    logic [8:0] PC_out;
    
// clock generation
    always #10 clk = ~ clk ;
    
// reset Generation
    initial begin
        clk = 0;
        reset = 1;
        #25 reset =0;
    end
    
    RISC_V tb_RISC_V (
        .clk(clk),
        .reset(reset),
        .ALU_Result(tb_ALU_Result),
        .INS_out(INS_out),
        .mux_out(mux_out),
        .rd1_out(rd1_out),
        .rd2_out(rd2_out),
        .PC_out(PC_out)
        );
        
    initial begin
        #2000;
        $finish ;
    end
endmodule
